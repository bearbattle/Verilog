module pipeline(
    input clk,
    input [31:0] A1,
    input [31:0] A2,
    input [31:0] B1,
    input [31:0] B2,
    output reg [31:0] C = 0);

endmodule
