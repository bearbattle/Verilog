`timescale 1ns / 1ps

module hazard(
    output reg [1:0] FALUAE,
    output reg [1:0] FALUBE
);



endmodule // hazard