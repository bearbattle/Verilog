`timescale 1ns / 1ps
module pc(
           input clk,
           input Reset,
           input [31:0] nPC,
           output reg [31:0] InstructionAddress
       );



endmodule // pc
