`timescale 1ns / 1ps

module alu(
    input A
);

endmodule // alu